module top_module(output zero);// Module body starts after semicolon
	assign zero = 0;
endmodule


assign one = 1'b1;
assign zero = 1'b0;

{3'b111, 3'b000} => 6'b111000
