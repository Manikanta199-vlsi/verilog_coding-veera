module top_module(output zero);// Module body starts after semicolon
	assign zero = 0;
endmodule


assign one = 1'b1;
